module tb_fake_n64_controller();
endmodule