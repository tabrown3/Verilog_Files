module tb_t_rex();

endmodule