module fake_n64_controller();
endmodule