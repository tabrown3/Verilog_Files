module filter_out_console_data(
    input data,
    input clk,
    output console_data
);

endmodule