module t_rex();

endmodule